library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MinhaPrimeiraAulaVHDL is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end MinhaPrimeiraAulaVHDL;

architecture rtl of MinhaPrimeiraAulaVHDL is

begin

end architecture;